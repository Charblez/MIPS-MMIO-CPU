// //----------------------------------------------------------------------------------------------------
// // Filename: SoC.sv
// // Author: Charles Bassani
// // Description: All components of chip connected
// //----------------------------------------------------------------------------------------------------
// `timescale 1ns/1ps

// //----------------------------------------------------------------------------------------------------
// // Module Declaration
// //----------------------------------------------------------------------------------------------------
// module SoC
// (

// );

// //----------------------------------------------------------------------------------------------------
// // Module Registers
// //----------------------------------------------------------------------------------------------------

// //----------------------------------------------------------------------------------------------------
// // Nested Modules
// //----------------------------------------------------------------------------------------------------
// DualChannelMem dpram_inst
// (
//     .clk(),
    
//     .we_a(),
//     .wdata_a(),
//     .rdata_a(),

//     .we_b(),
//     .wdata_b(),
//     .rdata_b()
// );

// //----------------------------------------------------------------------------------------------------
// // Module Logic
// //----------------------------------------------------------------------------------------------------
// endmodule